module hello();
    initial begin
        $display("hello from docker vivado");
        $finish;
    end
endmodule
